library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use ieee.std_logic_textio.all;

entity rom is
  port (
    ce       : in  std_logic;
    oe       : in  std_logic;
    byte_sel : in  std_logic_vector(3 downto 0);
    addr     : in  std_logic_vector(15 downto 0);
    data_out : out std_logic_vector(31 downto 0));
end entity rom;

architecture rtl of rom is

  type rom_bank_t is array (0 to 255) of std_logic_vector(31 downto 0);

  signal rom_bank_0 : rom_bank_t :=
    (
      "00000000001000100001100000100010",  -- SUB $r3, $r0, $r1	
      "00100000000000010000000000011001",  -- ADDI $r1, $r0, 24
      "00001000000000000000000000000010",  -- J to 0x0004 
      "10101010101010101010101010101010",  
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010",
      "10101010101010101010101010101010"
      );

begin  -- architecture rtl

  read : process (ce, oe, byte_sel, addr, rom_bank_0) is
  begin  -- process read
    if ce = '1' and oe = '1' then
      if byte_sel = "1111" then
        data_out <= rom_bank_0(to_integer(unsigned(addr(9 downto 2))));
      else
        data_out <= (others => '0');
      end if;
    else
      data_out <= (others => 'Z');
    end if;
  end process read;
end architecture rtl;
